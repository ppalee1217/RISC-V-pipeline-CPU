library verilog;
use verilog.vl_types.all;
entity compressor4_2_52 is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        d               : in     vl_logic;
        cin             : in     vl_logic;
        cout            : out    vl_logic;
        sum             : out    vl_logic;
        carry           : out    vl_logic
    );
end compressor4_2_52;
