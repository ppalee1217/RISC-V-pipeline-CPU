library verilog;
use verilog.vl_types.all;
entity blue_cell_19 is
    port(
        p2              : in     vl_logic;
        g1              : in     vl_logic;
        g2              : in     vl_logic;
        G               : out    vl_logic
    );
end blue_cell_19;
