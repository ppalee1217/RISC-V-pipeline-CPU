library verilog;
use verilog.vl_types.all;
entity black_cell_9 is
    port(
        p1              : in     vl_logic;
        p2              : in     vl_logic;
        g1              : in     vl_logic;
        g2              : in     vl_logic;
        G               : out    vl_logic;
        P               : out    vl_logic
    );
end black_cell_9;
